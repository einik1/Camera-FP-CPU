kobi_line_inst : kobi_line PORT MAP (
		clken	 => clken_sig,
		clock	 => clock_sig,
		shiftin	 => shiftin_sig,
		shiftout	 => shiftout_sig,
		taps0x	 => taps0x_sig,
		taps1x	 => taps1x_sig,
		taps2x	 => taps2x_sig,
		taps3x	 => taps3x_sig,
		taps4x	 => taps4x_sig
	);
